/*
 *      GEOFF MODULE
 *  (geometry_xy_plotter)
 *
<<<<<<< HEAD
 *       v 0.95. October 3rd, 2020
 * 
 * Geo-plotter/polyplot, sorter and blitter portions written by Brian Guralnick
 * Now inclused 12 bit fractional X&Y zoom and shrink scaling blitter operation.
=======
 *       v 0.1.001
>>>>>>> e95a3e278b115b0ea9f980c63d48b6bfbcc232d1
 *
 */

module geometry_xy_plotter (
<<<<<<< HEAD
    input wire clk,               // System clock
    input wire reset,             // Force reset
    input wire fifo_cmd_ready,    // 16-bit Data Command Ready signal
    input wire [15:0] fifo_cmd_in,// 16-bit Data Command bus
    input wire draw_busy,         // HIGH when pixel writer is busy, so geometry plotter will pause before sending any new pixels
    
    output wire load_cmd,         // HIGH when ready to receive next cmd_data[15:0] input
    output wire draw_cmd_rdy,     // Pulsed HIGH when data on draw_cmd[15:0] is ready to send to the pixel writer module
    output wire [35:0] draw_cmd,  // Bits [35:32] hold AUX function number 0-15:
=======
    input wire clk,              // System clock
    input wire reset,            // Force reset
    input wire fifo_cmd_ready,   // 16-bit Data Command Ready signal
    input wire [15:0] fifo_cmd_in,// 16-bit Data Command bus
    input wire draw_busy,        // HIGH when pixel writer is busy, so geometry plotter will pause before sending any new pixels
    
    output wire load_cmd,        // HIGH when ready to receive next cmd_data[15:0] input
    output wire draw_cmd_rdy,    // Pulsed HIGH when data on draw_cmd[15:0] is ready to send to the pixel writer module
    output wire [35:0] draw_cmd, // Bits [35:32] hold AUX function number 0-15:
    output wire fifo_cmd_busy    // HIGH when FIFO is full/nearly full
>>>>>>> e95a3e278b115b0ea9f980c63d48b6bfbcc232d1
    //  AUX=0  : Do nothing
    //  AUX=1  : Write pixel,                             : 31:24 color         : 23:12 Y coordinates : 11:0 X coordinates
    //  AUX=2  : Write pixel with color 0 mask,           : 31:24 color         : 23:12 Y coordinates : 11:0 X coordinates
    //  AUX=3  : Write from read pixel,                   : 31:24 ignored       : 23:12 Y coordinates : 11:0 X coordinates
    //  AUX=4  : Write from read pixel with color 0 mask, : 31:24 ignored       : 23:12 Y coordinates : 11:0 X coordinates
    //  AUX=6  : Read source pixel,                       : 31:24 ignored       : 23:12 Y coordinates : 11:0 X coordinates
    //  AUX=7  : Set Truecolor pixel color                : 31:24 8 bit alpha blend mix value : bits 23:0 hold RGB 24 bit color
<<<<<<< HEAD
    //                                                      Use function Aux3/4 to draw this color, only works if the destination is set to 16 bit true-color mode
=======
    //                                                    Use function Aux3/4 to draw this color, only works if the destination is set to 16 bit true-color mode
>>>>>>> e95a3e278b115b0ea9f980c63d48b6bfbcc232d1

    //  AUX=10 ; Resets the Write Pixel collision counter           : 31:24 sets transparent masked out color : bits 23:0 in true color mode, this holds RGB 24 bit mask color, in 8 bit mode, this allows for 3 additional transparent colors
    //  AUX=11 ; Resets the Write from read pixel collision counter : 31:24 sets transparent masked out color : bits 23:0 in true color mode, this holds RGB 24 bit mask color, in 8 bit mode, this allows for 3 additional transparent colors

    //  AUX=12 : Set destination raster width in bytes    : 15:0 holds destination raster image width in #bytes so the proper memory address can be calculated from the X&Y coordinates
    //  AUX=13 : Set source raster width in bytes,        : 15:0 holds source raster image width in #bytes so the proper memory address can be calculated from the X&Y coordinates
<<<<<<< HEAD
    //  AUX=14 : Set destination mem address,             : 31:24 bitplane mode : 23:0 hold destination base memory address for write pixel
    //  AUX=15 : Set source mem address,                  : 31:24 bitplane mode : 23:0 hold the source base memory address for read source pixel
    output wire fifo_cmd_busy     // HIGH when FIFO is full/nearly full
);

parameter int FIFO_MARGIN         = 32 ; // The number of extra commands the fifo has room after the 'fifo_cmd_busy' goes high
=======
    //  AUX=14 : Set destination mem address,             : 31:24 bitplane mode : 23:0 hold destination base memory addres for write pixel
    //  AUX=15 : Set source mem address,                  : 31:24 bitplane mode : 23:0 hold the source base memory address for read source pixel
);

parameter int FIFO_MARGIN         = 32 ; // The number of extra commadns the fifo has room after the 'fifo_cmd_busy' goes high
>>>>>>> e95a3e278b115b0ea9f980c63d48b6bfbcc232d1

logic [3:0] CMD_OUT_NOP           = 0  ;
logic [3:0] CMD_OUT_PXWRI         = 1  ;
logic [3:0] CMD_OUT_PXWRI_M       = 2  ;
logic [3:0] CMD_OUT_PXPASTE       = 3  ;
logic [3:0] CMD_OUT_PXPASTE_M     = 4  ;

logic [3:0] CMD_OUT_PXCOPY        = 6  ;
logic [3:0] CMD_OUT_SETARGB       = 7  ;

logic [3:0] CMD_OUT_RST_PXWRI_M   = 10 ;
logic [3:0] CMD_OUT_RST_PXPASTE_M = 11 ;
<<<<<<< HEAD

=======
>>>>>>> e95a3e278b115b0ea9f980c63d48b6bfbcc232d1
logic [3:0] CMD_OUT_DSTRWDTH      = 12 ;
logic [3:0] CMD_OUT_SRCRWDTH      = 13 ;
logic [3:0] CMD_OUT_DSTMADDR      = 14 ;
logic [3:0] CMD_OUT_SRCMADDR      = 15 ;

<<<<<<< HEAD
logic [7:0]  command_in     ;
logic [11:0] command_data12 ;
logic [7:0]  command_data8  ;

logic signed [11:0] x[0:3]      ; // 2-dimensional 12-bit register for x0-x3
logic signed [11:0] y[0:3]      ; // 2-dimensional 12-bit register for y0-y3
logic signed [11:0] max_x       ; // this reg will be both in this module and the memory pixel writer
logic signed [11:0] max_y       ; // this reg will be both in this module and the memory pixel writer

logic signed [23:0] blit_dest_x       ; // 
logic signed [11:0] blit_dest_x_int   ; // 
logic signed [23:0] blit_dest_rst_x   ; // 
logic signed [23:0] blit_dest_y       ; // 
logic signed [11:0] blit_dest_y_int   ; // 
logic signed [23:0] blit_dest_rst_y   ; // 
logic signed [23:0] blit_source_x     ; // 
logic signed [23:0] blit_source_y     ; // 
logic signed [11:0] blit_source_ofs_x ; // 
logic signed [11:0] blit_source_ofs_y ; // 
logic        [11:0] blit_width        ; // this stores how many pixels wide the blitter will copy
logic        [11:0] blit_height       ; // this stores how many pixels high the blitter will copy
logic               blit_running      ; // high when the blitter is running
logic               blit_paste_phase  ; // high when the blitter is running
logic signed [11:0] blit_dxs[0:3]     ; // Holds all the possible blitter starting paste X coordinates depending on selected paste features
logic signed [11:0] blit_dys[0:3]     ; // Holds all the possible blitter starting paste Y coordinates depending on selected paste features
logic        [12:0] blit_src_scale_x  ; // Holds the X blitter source upscale fraction, IE zoom ratio (4096:blit_src_scale_x), values 4095 through 1, or 4096 for off.
logic        [12:0] blit_src_scale_y  ; // Holds the Y blitter source upscale fraction, IE zoom ratio (4096:blit_src_scale_y), values 4095 through 1, or 4096 for off.
logic        [12:0] blit_dest_scale_x ; // Holds the X blitter destination downscale fraction, IE zoom ratio (blit_dest_scale_x:4096), values 4095 through 1, or 4096 for off.
logic        [12:0] blit_dest_scale_y ; // Holds the Y blitter destination downscale fraction, IE zoom ratio (blit_dest_scale_y:4096), values 4095 through 1, or 4096 for off.

logic [3:0]  draw_cmd_func        ;
logic [7:0]  draw_cmd_data_color  ;
logic [11:0] draw_cmd_data_word_Y ;
logic [11:0] draw_cmd_data_word_X ;
logic        draw_cmd_tx = 1'b0   ;

//************************************************************************************************************************************************
// Source command fifo
//************************************************************************************************************************************************
logic [15:0] cmd_data       ;
logic        fifo_cmd_rdy_n ;
=======
wire [7:0]  command_in     ;
wire [11:0] command_data12 ;
wire [7:0]  command_data8  ;

assign command_in     [7:0] = cmd_data[15:8] ;
assign command_data12[11:0] = cmd_data[11:0] ;
assign command_data8  [7:0] = cmd_data[7:0]  ;

reg [11:0] x[3:0] ; // 2-dimensional 12-bit register for x0-x3
reg [11:0] y[3:0] ; // 2-dimensional 12-bit register for y0-y3
reg [11:0] max_x  ; // this reg will be both in this module and the memory pixel writer
reg [11:0] max_y  ; // this reg will be both in this module and the memory pixel writer

reg [3:0]  draw_cmd_func        ;
reg [7:0]  draw_cmd_data_color  ;
reg [11:0] draw_cmd_data_word_Y ;
reg [11:0] draw_cmd_data_word_X ;
reg        draw_cmd_tx = 1'b0   ;

//************************************************
// Assign output port wires to internal registers
//************************************************
assign draw_cmd[35:32] = draw_cmd_func[3:0]         ;
assign draw_cmd[31:24] = draw_cmd_data_color[7:0]   ;
assign draw_cmd[23:12] = draw_cmd_data_word_Y[11:0] ;
assign draw_cmd[11:0]  = draw_cmd_data_word_X[11:0] ;
assign draw_cmd_rdy    = draw_cmd_tx && !draw_busy  ;

//************************************************
// geometry sequencer controls
//************************************************
reg [3:0]    geo_shape;            // 0 through 7 will draw their assigned shape, 8 through 15 will have different copy algorithms
reg          geo_fill;             // The geometric shape should be filled when set high
reg          geo_mask;             // If high, when drawing, the colors set in the 'collision counter' will not be drawn.
reg          geo_paste;            // If high, when drawing a geometric object, CMD_OUT_PXPASTE/_M will be used instead of CMD_OUT_PXWRI/_M for true color 16bit pixels
reg          geo_run   = 1'b0;     // High when a geometric shape is being drawn
reg [7:0]    geo_color;            // 8 bit pen drawing color

assign       load_cmd = ~geo_run;  // assigns the load_cmd output.  When the geometry unit is not drawing, the load_cmd goes high to load the next command.

//************************************************
// geometry counters
//************************************************
logic signed [11:0]   geo_x          ;
logic signed [11:0]   geo_y          ;
logic signed [11:0]   geo_xdir       ;
logic signed [11:0]   geo_ydir       ;
logic        [3:0]    geo_sub_func1  ; // auxiliary sequence counter
logic        [3:0]    geo_sub_func2  ; // auxiliary sequence counter
logic signed [11:0]   dx             ;
logic signed [11:0]   dy             ;
logic signed [11:0]   errd           ;
logic        [15:0]   cmd_data       ;
logic                 fifo_cmd_rdy_n ;
>>>>>>> e95a3e278b115b0ea9f980c63d48b6bfbcc232d1

scfifo  scfifo_component (
    .sclr        (reset),                                     // reset input
    .clock       (clk),                                       // system clock
<<<<<<< HEAD
    .wrreq       (fifo_cmd_ready),                            // connect this to the 'strobe' on the selected high.low Z80 bus output port
    .data        (fifo_cmd_in),                               // connect this to the 16 bit output port on the Z80 bus
    .almost_full (fifo_cmd_busy),                             // send to a selected bit on the Z80 status read port

    .empty       (fifo_cmd_rdy_n),                            // when LOW, the FIFO has commands for the geometry unit to process
    .rdreq       (load_cmd && !draw_busy),                    // connect to the listed inputs
    .q           (cmd_data[15:0]),                            // to geometry_xy_plotter cmd_data input
=======
    .wrreq       (fifo_cmd_ready),                            // connect this to the 'strobe' on the selected high.low Z80 bus output port.
    .data        (fifo_cmd_in),                               // connect this to the 16 bit output port on the Z80 bus.
    .almost_full (fifo_cmd_busy),                             // send to a selected bit on the Z80 status read port

    .empty       (fifo_cmd_rdy_n),                            // remember, when low, the FIFO has commands for the geometry unit to process
    .rdreq       (load_cmd && !draw_busy && !fifo_cmd_rdy_n), // connect to the listed inputs.
    .q           (cmd_data[15:0]),                            // to geometry_xy_plotter cmd_data input.
>>>>>>> e95a3e278b115b0ea9f980c63d48b6bfbcc232d1
    .full        ()                                           // optional, unused
);

defparam
    scfifo_component.add_ram_output_register = "ON",
    scfifo_component.almost_full_value       = (512 - FIFO_MARGIN),
    scfifo_component.intended_device_family  = "Cyclone IV",
    scfifo_component.lpm_hint                = "RAM_BLOCK_TYPE=M9K",
    scfifo_component.lpm_numwords            = 512,
    scfifo_component.lpm_showahead           = "ON",
    scfifo_component.lpm_type                = "scfifo",
    scfifo_component.lpm_width               = 16,
    scfifo_component.lpm_widthu              = 9,
    scfifo_component.overflow_checking       = "ON",
    scfifo_component.underflow_checking      = "ON",
    scfifo_component.use_eab                 = "ON";

<<<<<<< HEAD
//************************************************************************************************************************************************
// Source command coordinate sorting and interpretation pipe.
//************************************************************************************************************************************************
logic                sort_cmd_rdy      ;
logic [15:0]         sort_data_pipe    ; // cmd_data pipeline OUT from poly_sort into geo_xy_plotter
logic signed  [11:0] sort_coords[0:15] ; // array package of sorted coordinates for the linegen
logic signed  [11:0] sort_y_range[0:1] ; // array package of defining the starting and ending Y coordinates for a filled polygon
logic [1:0]          lg_seq_size[0:1]  ;
logic                lg_fill           ;
logic                draw_shape        ;
logic [7:0]          blit_features     ;
logic [7:0]          blit_mask_col     ;


//************************************************************************************************************************************************
// Geometry XY line plotter.
//************************************************************************************************************************************************
logic                plot_cmd_rdy       ;
logic [15:0]         plot_data_pipe     ; // cmd_data pipeline OUT from poly_plot into the blitter
logic signed  [11:0] plot_pixel_xy[0:1] ; // xy coordinates to plot to
logic                plot_pixel_ena     ;
logic [7:0]          plot_pixel_col     ;
logic                plot_busy          ;
logic [7:0]          p_blit_features    ;
logic [7:0]          p_blit_mask_col    ;

poly_plot plotter (
// inputs
    .clk               ( clk             ),
    .reset             ( reset           ),
    .enable            ( !draw_busy      ), // !pixel_writer busy input
    .blitter_busy      ( blit_running    ),
    .cmd_rdy_in        ( !fifo_cmd_rdy_n ),
    .cmd_in            ( cmd_data        ), // ** cmd_data pipeline input from FIFO
    .x_in              ( x               ), // xy[0,1,2,3] registers
    .y_in              ( y               ), // xy[0,1,2,3] registers
//outputs
    .pixel_ena         ( plot_pixel_ena  ),
    .pixel_xy          ( plot_pixel_xy   ),  // array package of sorted coordinates for the linegen 0&1
    .pixel_col         ( plot_pixel_col  ),  // array package of sorted coordinates for the linegen 0&1
    .plotter_busy      ( plot_busy       ),  // array containing the number of line coordinates for each linegen to run
    .blit_features_out ( p_blit_features ),  // Tells the blitter module to copy & paste a rectangle.
    .blit_mask_col_out ( p_blit_mask_col ),  // Tells the blitter copy pixel function how to transpose the source pixel color
    .blit_src_scale_x  ( blit_src_scale_x),  // Holds the X blitter source upscale fraction, IE zoom ratio (4096:blit_src_scale_x), values 4095 through 1, or 4096 for off.
    .blit_src_scale_y  ( blit_src_scale_y),  // Holds the Y blitter source upscale fraction, IE zoom ratio (4096:blit_src_scale_y), values 4095 through 1, or 4096 for off.
    .blit_dest_scale_x ( blit_dest_scale_x), // Holds the X blitter destination downscale fraction, IE zoom ratio (blit_dest_scale_x:4096), values 4095 through 1, or 4096 for off.
    .blit_dest_scale_y ( blit_dest_scale_y)  // Holds the Y blitter destination downscale fraction, IE zoom ratio (blit_dest_scale_y:4096), values 4095 through 1, or 4096 for off.
);


//************************************************************************************************************************************************
// Geometry plotter address & pointers command decoder and registers,
// final pixel blitter & command output to address generator.
//************************************************************************************************************************************************

always_comb begin

    // Assign output port wires to internal registers
    draw_cmd[35:32]      = draw_cmd_func[3:0]         ;
    draw_cmd[31:24]      = draw_cmd_data_color[7:0]   ;
    draw_cmd[23:12]      = draw_cmd_data_word_Y[11:0] ;
    draw_cmd[11:0]       = draw_cmd_data_word_X[11:0] ;
    draw_cmd_rdy         = draw_cmd_tx && !draw_busy  ;

    // Break out cmd_data bus into logical words
    command_in     [7:0] = cmd_data[15:8]        ;
    command_data12[11:0] = cmd_data[11:0]        ;
    command_data8  [7:0] = cmd_data[7:0]         ;

    // Assign the load_cmd output - when the geometry unit is not drawing, the load_cmd goes high to load the next command
    load_cmd             = !plot_busy  && !fifo_cmd_rdy_n  && !blit_running ;

// Setup all the possible blitter starting X&Y coordinates based on which feature are enabled
blit_dxs[3] = plot_pixel_xy[0]+blit_width[10:1]  ; // Beginning paste X coordinates with Mirror enabled  and Center Paste enabled
blit_dxs[2] = plot_pixel_xy[0]+blit_width[10:0]  ; // Beginning paste X coordinates with Mirror enabled  and Center Paste disabled
blit_dxs[1] = plot_pixel_xy[0]-blit_width[10:1]  ; // Beginning paste X coordinates with Mirror disabled and Center Paste enabled
blit_dxs[0] = plot_pixel_xy[0]                   ; // Beginning paste X coordinates with Mirror disabled and Center Paste disabled

blit_dys[3] = plot_pixel_xy[1]+blit_height[10:1] ; // Beginning paste Y coordinates with Flip enabled  and Center Paste enabled
blit_dys[2] = plot_pixel_xy[1]+blit_height[10:0] ; // Beginning paste Y coordinates with Flip enabled  and Center Paste disabled
blit_dys[1] = plot_pixel_xy[1]-blit_height[10:1] ; // Beginning paste Y coordinates with Flip disabled and Center Paste enabled
blit_dys[0] = plot_pixel_xy[1]                   ; // Beginning paste Y coordinates with Flip disabled and Center Paste disabled

// Assign integer only versions of the destination coordinates for the blitter paste coordinates.
blit_dest_x_int = blit_dest_x[23:12];
blit_dest_y_int = blit_dest_y[23:12];

end // always_comb

always_ff @(posedge clk or posedge reset) begin
=======
logic linegen_start       ;
logic line_done           ;
logic pass_thru_a         ;
logic pass_thru_b         ;
logic y_stop              ;
logic y_stopped           ;
logic [11:0] y_stop_coord ;
logic line_dat_rdy        ;
logic line_gen_running    ;
logic [11:0] gen_x        ;
logic [11:0] gen_y        ;

line_generator linegen_1 (
// inputs
  .clk            ( clk ),              // 125 MHz pixel clock
  .reset          ( reset ),            // asynchronous reset
  .run            ( linegen_start ),    // HIGH during drawing
  .draw_busy      ( draw_busy ),        // draw_busy input from parent module
  .pass_thru_a    ( pass_thru_a ),      // set HIGH to pass through aX/aY coordinates
  .pass_thru_b    ( pass_thru_b ),      // set HIGH to pass through bX/bY coordinates
  .aX             ( x[0] ),             // 12-bit X-coordinate for line start
  .aY             ( y[0] ),             // 12-bit Y-coordinate for line start
  .bX             ( x[1] ),             // 12-bit X-coordinate for line end
  .bY             ( y[1] ),             // 12-bit Y-coordinate for line end
  .ena_stop_y     ( y_stop ),           // set HIGH to make line generator stop at stop_ypos
  .stop_ypos      ( y_stop_coord ),     // Y_coordinate to stop at
// outputs
  .busy           ( line_gen_running ), // HIGH when line_generator is running
  .X_coord        ( gen_x ), // 12-bit X-coordinate for current pixel
  .Y_coord        ( gen_y ), // 12-bit Y-coordinate for current pixel
  .pixel_data_rdy ( line_dat_rdy ),     // HIGH when coordinate outputs are valid
  .ypos_stopped   ( y_stopped ),        // HIGH when stopped on Y-position
  .line_complete  ( line_done )         // HIGH when line is completed

);

always @(posedge clk or posedge reset) begin
>>>>>>> e95a3e278b115b0ea9f980c63d48b6bfbcc232d1

    if (reset) begin    // reset to defaults
        
        // reset coordinate registers
        for ( integer i = 0; i < 4; i++ ) begin
<<<<<<< HEAD
            x[i] <= { 12'b0 } ;
            y[i] <= { 12'b0 } ;
        end
        
        max_x                <= 12'b0 ;
        max_y                <= 12'b0 ;
        
        blit_dest_x         <= 12'b0 ; // 
        blit_dest_rst_x     <= 12'b0 ; // 
        blit_dest_y         <= 12'b0 ; // 
        blit_source_x       <= 12'b0 ; // 
        blit_source_y       <= 12'b0 ; // 
        blit_source_ofs_x   <= 12'b0 ; // 
        blit_source_ofs_y   <= 12'b0 ; // 
        blit_width          <= 12'b0 ; // this stores how many pixels wide the blitter will copy
        blit_height         <= 12'b0 ; // this stores how many pixels high the blitter will copy
        blit_running        <= 1'b0 ;  // high when the blitter is running
        blit_paste_phase    <= 1'b0 ;  // high when the blitter is pasting, low when copying
=======
            x[i]  <= { 12'b0 } ;
            y[i]  <= { 12'b0 } ;
        end
        max_x     <= 12'b0     ;
        max_y     <= 12'b0     ;
>>>>>>> e95a3e278b115b0ea9f980c63d48b6bfbcc232d1

        // reset draw command registers
        draw_cmd_func        <= 4'b0  ;
        draw_cmd_data_color  <= 8'b0  ;
        draw_cmd_data_word_Y <= 12'b0 ;
        draw_cmd_data_word_X <= 12'b0 ;
        draw_cmd_tx          <= 1'b0  ;
<<<<<<< HEAD
        
        
    end else if (!draw_busy) begin  // Everything must PAUSE if the incoming draw_busy signal from the pixel_writer is high
     
        
//************************************************************************************************************************************************
// When the plotter is busy, pass the output coordinates as a draw command.
// If the blitter is enables, use the plot coordinates as the center of a COPY, the PASTE command
// sequence with a box size of blit_width & blit_height.
//************************************************************************************************************************************************
   if (plot_busy || blit_running ) begin

//************************************************************************************************************************************************
// p_blit_features bitmask features:
// 0 = Enable blitter         1 = run biltter copying source to output coordinates, 0 = Simple pixel write command
// 1 = Enable paste mask      1 = Paste pixels with transparency mask, 0 = Always paste pixels even if the source pixel is the selected transparent color
// 2 = Enable H-center paste  1 = Offset the paste to the left by half of blit_width, 0 = Use the paste coordinates as the left margin
// 3 = Enable Mirror paste    1 = Mirror the output on the X axis.
// 4 = Enable V-center paste  1 = Offset the paste up by half of blit_height, 0 = Use the paste coordinates as the first line of the paste
// 5 = Enable Flip paste      1 = Flip the output on the Y axis.
// 6 = Enable Rotate 90 degree paste  1 = Swaps the X&Y coordinates on the paste.
// 7 = Enable Rotate 45 degree paste  1 = Increments/decrements the X&Y coordinates on the paste in unison.
//************************************************************************************************************************************************
if ( !p_blit_features[0] ) begin // ***** Blitter disabled.
        if ( plot_pixel_ena && ( plot_pixel_xy[0] >= 0 && plot_pixel_xy[0] < max_x ) && ( plot_pixel_xy[1] >=0 && plot_pixel_xy[1] < max_y ) ) begin
            blit_running         <= 1'b0;
            draw_cmd_func        <= CMD_OUT_PXWRI    ;
            draw_cmd_data_word_X <= plot_pixel_xy[0] ; // ... at X-coordinate
            draw_cmd_data_word_Y <= plot_pixel_xy[1] ; // ... and Y-coordinate
            draw_cmd_data_color  <= plot_pixel_col   ;    
            draw_cmd_tx          <= 1'b1             ; // let PAGET know valid pixel data is incoming
        end
        else draw_cmd_tx         <= 1'b0 ; // otherwise turn off draw command

end else begin // ***** Blitter enabled.

        if (!blit_running && plot_pixel_ena ) begin   // Blitter isn't yet running, so, initialize it.
            blit_running         <= 1'b1  ;           // Signal blitter running so the poly_plot module knows to wait for the copy/paste.
            blit_source_x        <= 24'd0 ;           // Clear the source coordinates
            blit_source_y        <= 24'd0 ;
            blit_paste_phase     <= 1'b0  ;           // Tells the blitter that a copy pixel has been done and ready for a paste pixel

            // Set the initial destination coordinates based on the Enable center H/V, and mirror/flip blitter features.
            blit_dest_x[23:12]     <= blit_dxs[p_blit_features[3:2]] ; // Set the beginning paste X coordinates.
            blit_dest_rst_x[23:12] <= blit_dxs[p_blit_features[3:2]] ; // tells the copy where to reset X during a Y increment
            blit_dest_y[23:12]     <= blit_dys[p_blit_features[5:4]] ; // Set the beginning paste Y coordinates.
            blit_dest_rst_y[23:12] <= blit_dys[p_blit_features[5:4]] ; // tells the copy where to reset Y during a X increment when copying with a 90 degree rotation
            // clear the floating point locations
            blit_dest_x[11:0]      <= 12'd0                          ; // Set the beginning paste X coordinates.
            blit_dest_rst_x[11:0]  <= 12'd0                          ; // tells the copy where to reset X during a Y increment
            blit_dest_y[11:0]      <= 12'd0                          ; // Set the beginning paste Y coordinates.
            blit_dest_rst_y[11:0]  <= 12'd0                          ; // tells the copy where to reset Y during a X increment when copying with a 90 degree rotation
            
         end else if ( blit_running ) begin // Blitter has been setup, now in running mode

         //  Whether reading or writing a pixel, if the destination pixel is inside the valid screen coordinates, enable the draw command TX
            if ( (blit_dest_x_int >= 0 && blit_dest_x_int < max_x ) && ( blit_dest_y_int >=0 && blit_dest_y_int < max_y ) ) draw_cmd_tx <= 1'b1 ;
         //  Otherwise stop the draw command TX
            else                                                                                                            draw_cmd_tx <= 1'b0 ;

         // During the first blitter phase, set the output command to the copy pixel coordinates and set the next phase to a paste pixel
                        if (!blit_paste_phase) begin
                        draw_cmd_func        <= CMD_OUT_PXCOPY   ;                         // Copy the source pixel command.
                        draw_cmd_data_word_X <= blit_source_x[23:12] + blit_source_ofs_x ; // ... at X-coordinate
                        draw_cmd_data_word_Y <= blit_source_y[23:12] + blit_source_ofs_y ; // ... and Y-coordinate
                        draw_cmd_data_color  <= p_blit_mask_col  ;                         // Copy color pixel transformation  (Read pixel is XORed with this number)   
                        blit_paste_phase     <= 1'b1 ;                                     // signal the next blitter phase, paste the copied pixel
                        end
            
         // During the second blitter phase, (PART 1) set the output command to the paste pixel coordinates.
                        if ( blit_paste_phase) begin
                        draw_cmd_func        <= p_blit_features[1] ? CMD_OUT_PXPASTE_M : CMD_OUT_PXPASTE ; // Write the pixel with the optional paste mask feature
                        draw_cmd_data_word_X <= blit_dest_x_int    ;                                       // ... at X-coordinate
                        draw_cmd_data_word_Y <= blit_dest_y_int    ;                                       // ... and Y-coordinate
                        draw_cmd_data_color  <= plot_pixel_col     ;                                       // Second XORed color transformation   
                        draw_cmd_tx          <= 1'b1               ;                                       // let PAGET know valid pixel data is incoming
                        end

         // During the second blitter phase, (PART 2), OR when the destination paste pixel coordinates are OUTSIDE the valid screen coordinates,
         // (this step skipps a clock cycle when addressing pixels off the screen area)
         // Increment/decrement all the X&Y pointers/coordinates and set the blitter phase back into copy pixel mode.
         
         if ( blit_paste_phase || !( (blit_dest_x_int >= 0 && blit_dest_x_int < max_x ) && ( blit_dest_y_int >=0 && blit_dest_y_int < max_y ) ) ) begin

              blit_paste_phase     <= 1'b0 ;  // signal the next blitter phase, copy pixel.
         
                        if ( blit_source_x[23:12] == blit_width && blit_source_y[23:12] == blit_height ) begin // the copy has reached the blit_width/height
                        blit_running         <= 1'b0            ; // turn off blitter
                        end else if ( blit_source_x[23:12] != blit_width ) begin // width has not been reached, increment the X coordinates
                                                           blit_source_x <= blit_source_x + blit_src_scale_x ;

                                                      if ( p_blit_features[7]) begin   // Paste with 45 degree rotate begin
                                                           if ( !p_blit_features[3] ) blit_dest_x   <= blit_dest_x + blit_dest_scale_x ; // Horizontal mirror off
                                                           else                       blit_dest_x   <= blit_dest_x - blit_dest_scale_x ; // Horizontal mirror on
                                                           if ( !p_blit_features[5] ) blit_dest_y   <= blit_dest_y + blit_dest_scale_y ; // Vertical flip off
                                                           else                       blit_dest_y   <= blit_dest_y - blit_dest_scale_y ; // Vertical flip on

                                                      end else begin                   // no Paste 45 degree rotate begin
                                                      if (!p_blit_features[6]) begin   // Paste un-rotated
                                                           if ( !p_blit_features[3] ) blit_dest_x   <= blit_dest_x + blit_dest_scale_x ; // Horizontal mirror off
                                                           else                       blit_dest_x   <= blit_dest_x - blit_dest_scale_x ; // Horizontal mirror on
                                                      end else begin                   // Paste rotated 90 degrees
                                                           if ( !p_blit_features[5] ) blit_dest_y   <= blit_dest_y + blit_dest_scale_y ; // Vertical flip off
                                                           else                       blit_dest_y   <= blit_dest_y - blit_dest_scale_y ; // Vertical flip on
                                                      end
                                                      end  //  no Paste 45 degree rotate end

                        end else begin // width has been reached, increment the Y coordinates and reset the X coordinates
                                                           blit_source_y <= blit_source_y + blit_src_scale_y ;

                                                      if ( p_blit_features[7]) begin  // Paste with 45 degree rotate
                                                           if ( !p_blit_features[5] ) blit_dest_y     <= blit_dest_rst_y + blit_dest_scale_y ; // Vertical flip off
                                                           else                       blit_dest_y     <= blit_dest_rst_y - blit_dest_scale_y ; // Vertical flip on
                                                           if ( !p_blit_features[5] ) blit_dest_x     <= blit_dest_rst_x - blit_dest_scale_x ; // New line return 
                                                           else                       blit_dest_x     <= blit_dest_rst_x + blit_dest_scale_x ; // New line return 
                                                           
                                                           if ( !p_blit_features[5] ) blit_dest_rst_x <= blit_dest_rst_x - blit_dest_scale_x ; // Modify new line return position 
                                                           else                       blit_dest_rst_x <= blit_dest_rst_x + blit_dest_scale_x ; // Modify new line return position 
                                                             
                                                           if ( !p_blit_features[3] ) blit_dest_x     <= blit_dest_rst_x - blit_dest_scale_x ; // Horizontal mirror off
                                                           else                       blit_dest_x     <= blit_dest_rst_x + blit_dest_scale_x ; // Horizontal mirror on
                                                           if ( !p_blit_features[3] ) blit_dest_y     <= blit_dest_rst_y + blit_dest_scale_y ; // New line return 
                                                           else                       blit_dest_y     <= blit_dest_rst_y - blit_dest_scale_y ; // New line return 
                                                           
                                                           if ( !p_blit_features[3] ) blit_dest_rst_y <= blit_dest_rst_y + blit_dest_scale_y ; // Modify new line return position 
                                                           else                       blit_dest_rst_y <= blit_dest_rst_y - blit_dest_scale_y ; // Modify new line return position 
                                                      
                                                      end else begin                   // Paste horizontal or vertical
                                                      if (!p_blit_features[6]) begin   // Paste un-rotated
                                                           if ( !p_blit_features[5] ) blit_dest_y   <= blit_dest_y + blit_dest_scale_y ; // Vertical flip off
                                                           else                       blit_dest_y   <= blit_dest_y - blit_dest_scale_y ; // Vertical flip on
                                                                                      blit_dest_x   <= blit_dest_rst_x                 ; // New line return  
                                                      end else begin                   // Paste rotated 90 degrees
                                                           if ( !p_blit_features[3] ) blit_dest_x   <= blit_dest_x + blit_dest_scale_x ; // Horizontal mirror off
                                                           else                       blit_dest_x   <= blit_dest_x - blit_dest_scale_x ; // Horizontal mirror on
                                                                                      blit_dest_y   <= blit_dest_rst_y                 ; // New line return  
                                                      end
                                                      end  //  no Paste 45 degree rotate end

                                                           blit_source_x <= 24'd0 ;
                        end
                        
            end // end of paste pixel phase
         end else draw_cmd_tx  <= 1'b0 ; // end of blitter running
     end // end of p_blit_features[0] enable

end else begin // end of plot_busy

        // This code interprets the incoming commands when the linegens and blitter are not generating pixels
        if ( load_cmd ) begin  // when the cmd_rdy input is LOW and the geometry unit geo_run is not running, execute the following command input
         
            casez (command_in)
             
                8'b10?????? : x[command_in[5:4]] <= command_data12 ;
                
                8'b11?????? : y[command_in[5:4]] <= command_data12 ;
                
                8'b011111?? : begin // set 24-bit destination screen memory pointer for plotting
                    draw_cmd_func        <= CMD_OUT_DSTMADDR[3:0]  ; // sets the output function
                    draw_cmd_data_color  <= command_data8          ; // set screen_mode (bits per pixel)
                    draw_cmd_data_word_Y <= y[command_in[1:0]]     ; // sets the upper 12 bits of the destination address
                    draw_cmd_data_word_X <= x[command_in[1:0]]     ; // sets the lower 12 bits of the destination address
                    draw_cmd_tx          <= 1'b1                   ; // transmits the command
                end
             
                8'b011110?? : begin // set 24-bit source screen memory pointer for blitter copy
                    draw_cmd_func        <= CMD_OUT_SRCMADDR[3:0]  ; // sets the output function
                    draw_cmd_data_color  <= command_data8          ; // set screen_mode (bits per pixel)
                    draw_cmd_data_word_Y <= y[command_in[1:0]]     ; // sets the upper 12 bits of the destination address
                    draw_cmd_data_word_X <= x[command_in[1:0]]     ; // sets the lower 12 bits of the destination address
                    draw_cmd_tx          <= 1'b1                   ; // transmits the command
                end
                
                 8'b0111011? : begin  // Sets the blitter source offset X&Y position with x/y[2&3]
                    blit_source_ofs_x    <= x[{1'b1,command_in[0]}]     ; // sets the upper 12 bits of the destination address
                    blit_source_ofs_y    <= y[{1'b1,command_in[0]}]     ; // sets the lower 12 bits of the destination address
                end

                 8'b0111010? : begin  // Sets the blitter copy width and height with x/y[2&3]
                    blit_width           <= x[{1'b1,command_in[0]}]     ; // sets the upper 12 bits of the destination address
                    blit_height          <= y[{1'b1,command_in[0]}]     ; // sets the lower 12 bits of the destination address
                end
              
                8'd115 : begin  // set the number of bytes per horizontal line in the destination raster
                    draw_cmd_func        <= CMD_OUT_DSTRWDTH[3:0]  ; // sets the output function
                    draw_cmd_data_color  <= command_data8          ; // set bitplane mode (bits per pixel)
                    draw_cmd_data_word_Y <= y[2]                   ; // null
                    draw_cmd_data_word_X <= x[2]                   ; // sets the lower 12 bits of the destination address
                    draw_cmd_tx          <= 1'b1                   ; // transmits the command
                end
                
                8'd114 : begin  // set the number of bytes per horizontal line in the source raster
                    draw_cmd_func        <= CMD_OUT_SRCRWDTH[3:0]  ; // sets the output function
                    draw_cmd_data_color  <= command_data8          ; // set bitplane mode (bits per pixel)
                    draw_cmd_data_word_Y <= y[2]                   ; // sets the lower 12 bits of the destination address
                    draw_cmd_data_word_X <= x[2]                   ; // null
                    draw_cmd_tx          <= 1'b1                   ; // transmits the command
                end
                    
                8'd113 : begin  // set the number of bytes per horizontal line in the destination raster
                    draw_cmd_func        <= CMD_OUT_DSTRWDTH[3:0]  ; // sets the output function
                    draw_cmd_data_color  <= command_data8          ; // set bitplane mode (bits per pixel)
                    draw_cmd_data_word_Y <= y[3]                   ; // null
                    draw_cmd_data_word_X <= x[3]                   ; // sets the lower 12 bits of the destination address
                    draw_cmd_tx          <= 1'b1                   ; // transmits the command
                end
                    
                8'd112 : begin  // set the number of bytes per horizontal line in the source raster
                    draw_cmd_func        <= CMD_OUT_SRCRWDTH[3:0]  ; // sets the output function
                    draw_cmd_data_color  <= command_data8          ; // set bitplane mode (bits per pixel)
                    draw_cmd_data_word_Y <= y[3]                   ; // sets the lower 12 bits of the destination address
                    draw_cmd_data_word_X <= x[3]                   ; // null
                    draw_cmd_tx          <= 1'b1                   ; // transmits the command
                end

                8'd95  : begin
                    max_x <= x[0] ;    // set max width & height of screen to x0/y0
                    max_y <= y[0] ;
=======

        // reset geometry sequencer controls
        geo_shape     <= 4'b0  ;
        geo_fill      <= 1'b0  ;
        geo_mask      <= 1'b0  ;
        geo_paste     <= 1'b0  ;
        geo_run       <= 1'b0  ;
        geo_color     <= 8'b0  ;
        linegen_start <= 1'b0  ;
        
        // reset geometry counters
        geo_x         <= 12'b0 ;
        geo_y         <= 12'b0 ;
        geo_xdir      <= 12'b0 ;
        geo_ydir      <= 12'b0 ;
        geo_sub_func1 <= 4'b0  ;
        geo_sub_func2 <= 4'b0  ;
        dx            <= 12'b0 ;
        dy            <= 12'b0 ;
        errd          <= 12'b0 ;

    end else if (!draw_busy) begin
    
        if ( !fifo_cmd_rdy_n && ~geo_run ) begin  // when the fifo_cmd_rdy_n input is LOW and the geometry unit geo_run is not running, execute the following command input

            casez (command_in)
            
                8'b10?????? : x[command_in[5:4]] <= command_data12;
                
                8'b11?????? : y[command_in[5:4]] <= command_data12;

                8'b011111?? : begin // set 24-bit destination screen memory pointer for plotting
                    draw_cmd_func        <= CMD_OUT_DSTMADDR[3:0];   // sets the output function
                    draw_cmd_data_color  <= command_data8;           // set screen_mode (bits per pixel)
                    draw_cmd_data_word_Y <= y[command_in[1:0]];      // sets the upper 12 bits of the destination address
                    draw_cmd_data_word_X <= x[command_in[1:0]];      // sets the lower 12 bits of the destination address
                    draw_cmd_tx          <= 1'b1;                    // transmits the command
                end

                8'b011110?? : begin // set 24-bit source screen memory pointer for blitter copy
                    draw_cmd_func        <= CMD_OUT_SRCMADDR[3:0];   // sets the output function
                    draw_cmd_data_color  <= command_data8;           // set screen_mode (bits per pixel)
                    draw_cmd_data_word_Y <= y[command_in[1:0]];      // sets the upper 12 bits of the destination address
                    draw_cmd_data_word_X <= x[command_in[1:0]];      // sets the lower 12 bits of the destination address
                    draw_cmd_tx          <= 1'b1;                    // transmits the command
                end
                    
                8'd119 : begin  //Ignore for now
                    //destmem <= x[11:0][0] * 4096 + y[11:0][0];  // set both source & destination pointers for blitter copy
                    //srcmem  <= x[11:0][1] * 4096 + y[11:0][1];
                end
                
                8'd118 : begin //Ignore for now
                    //destmem <= x[11:0][1] * 4096 + y[11:0][1];  // set both source & destination pointers for blitter copy
                    //srcmem  <= x[11:0][0] * 4096 + y[11:0][0];
                end
                
                8'd117 : begin //Ignore for now
                    //destmem <= x[11:0][2] * 4096 + y[11:0][2];  // set both source & destination pointers for blitter copy
                    //srcmem  <= x[11:0][3] * 4096 + y[11:0][3];
                end
                
                8'd116 : begin //Ignore for now
                    //destmem <= x[11:0][3] * 4096 + y[11:0][3];  // set both source & destination pointers for blitter copy
                    //srcmem  <= x[11:0][2] * 4096 + y[11:0][2];
                end
                        
                8'd115 : begin  // set the number of bytes per horizontal line in the destination raster
                    draw_cmd_func        <= CMD_OUT_DSTRWDTH[3:0];   // sets the output function
                    draw_cmd_data_color  <= command_data8;           // set bitplane mode (bits per pixel)
                    draw_cmd_data_word_Y <= y[2];                    // null
                    draw_cmd_data_word_X <= x[2];                    // sets the lower 12 bits of the destination address
                    draw_cmd_tx          <= 1'b1;                    // transmits the command
                end
                    
                8'd114 : begin  // set the number of bytes per horizontal line in the source raster
                    draw_cmd_func        <= CMD_OUT_SRCRWDTH[3:0];   // sets the output function
                    draw_cmd_data_color  <= command_data8;           // set bitplane mode (bits per pixel)
                    draw_cmd_data_word_Y <= y[2];                    // sets the lower 12 bits of the destination address
                    draw_cmd_data_word_X <= x[2];                    // null
                    draw_cmd_tx          <= 1'b1;                    // transmits the command
                end
                    
                8'd113 : begin  // set the number of bytes per horizontal line in the destination raster
                    draw_cmd_func        <= CMD_OUT_DSTRWDTH[3:0];   // sets the output function
                    draw_cmd_data_color  <= command_data8;           // set bitplane mode (bits per pixel)
                    draw_cmd_data_word_Y <= y[3];                    // null
                    draw_cmd_data_word_X <= x[3];                    // sets the lower 12 bits of the destination address
                    draw_cmd_tx          <= 1'b1;                    // transmits the command
                end
                    
                8'd112 : begin  // set the number of bytes per horizontal line in the source raster
                    draw_cmd_func        <= CMD_OUT_SRCRWDTH[3:0];   // sets the output function
                    draw_cmd_data_color  <= command_data8;           // set bitplane mode (bits per pixel)
                    draw_cmd_data_word_Y <= y[3];                    // sets the lower 12 bits of the destination address
                    draw_cmd_data_word_X <= x[3];                    // null
                    draw_cmd_tx          <= 1'b1;                    // transmits the command
                end

                    
                8'd95  : begin
                    max_x <= x[0];    // set max width & height of screen to x0/y0
                    max_y <= y[0];
>>>>>>> e95a3e278b115b0ea9f980c63d48b6bfbcc232d1
                    //********************  no command to be set......draw_cmd_tx <= 1'b1;
                end
                
                8'd94  : begin
<<<<<<< HEAD
                    max_x <= x[1] ;    // set max width & height of screen to x1/y1
                    max_y <= y[1] ;
=======
                    max_x <= x[1];    // set max width & height of screen to x1/y1
                    max_y <= y[1];
>>>>>>> e95a3e278b115b0ea9f980c63d48b6bfbcc232d1
                    //********************  no command to be set......draw_cmd_tx <= 1'b1;
                end
                
                8'd93  : begin
<<<<<<< HEAD
                    max_x <= x[2] ; // set max width & height of screen to x2/y2
                    max_y <= y[2] ;
=======
                    max_x <= x[2];    // set max width & height of screen to x2/y2
                    max_y <= y[2];
>>>>>>> e95a3e278b115b0ea9f980c63d48b6bfbcc232d1
                    //********************  no command to be set......draw_cmd_tx <= 1'b1;
                end
                
                8'd92 : begin
<<<<<<< HEAD
                    max_x <= x[3] ; // set max width & height of screen to x3/y3
                    max_y <= y[3] ;
=======
                    max_x <= x[3];    // set max width & height of screen to x3/y3
                    max_y <= y[3];
>>>>>>> e95a3e278b115b0ea9f980c63d48b6bfbcc232d1
                    //********************  no command to be set......draw_cmd_tx <= 1'b1;
                end
                        
                8'd91 : begin               // clear the pixel collision counter and sets all 3 transparent mask colors to 1 8-bit color in the source function data
<<<<<<< HEAD
                    draw_cmd_func        <= CMD_OUT_RST_PXWRI_M[3:0]                   ; // sets the output funtion
                    draw_cmd_data_color  <= command_data8                              ; // sets the mask color
                    draw_cmd_data_word_Y <= { command_data8[7:0], command_data8[7:4] } ; // sets mask color #2 and 1/2 or #3
                    draw_cmd_data_word_X <= { command_data8[3:0], command_data8[7:4] } ; // sets mask color 1/2 or #3 and #4
                    draw_cmd_tx          <= 1'b1                                       ; // transmits the command
                end
                
                8'd90 : begin               // clear the blitter copy pixel collision counter
                    draw_cmd_func        <= CMD_OUT_RST_PXPASTE_M[3:0]                 ; // sets the output funtion
                    draw_cmd_data_color  <= command_data8                              ; // sets the mask color
                    draw_cmd_data_word_Y <= { command_data8[7:0], command_data8[7:4] } ; // sets mask color #2 and 1/2 or #3
                    draw_cmd_data_word_X <= { command_data8[3:0], command_data8[7:4] } ; // sets mask color 1/2 or #3 and #4
                    draw_cmd_tx          <= 1'b1                                       ; // transmits the command
                end

                default : begin
                    draw_cmd_tx          <= 1'b0  ; // no command to transmit
                end

            endcase
            
        end else draw_cmd_tx          <= 1'b0  ; // !load_cmd
      end // !plot_busy
    end // !draw_busy

end //always @(posedge clk)

endmodule



/*
 * poly_plot module
 *
 * renders lines and fills
 *
 */
module poly_plot (
// inputs
    input logic                 clk              ,
    input logic                 reset            ,
    input logic                 enable           , // !pixel_writer busy input
    input logic                 blitter_busy     , // When high, pause the linegens
    input logic                 cmd_rdy_in       ,
    input logic          [15:0] cmd_in           ,
    input logic   signed [11:0] x_in [0:3]       , // values to plot
    input logic   signed [11:0] y_in [0:3]       , // values to plot
//outputs
    output logic                pixel_ena        ,
    output logic         [7:0]  pixel_col        ,
    output logic  signed [11:0] pixel_xy [0:1]   , // Destination coordinates
    output logic                plotter_busy     , // The linegens are running
    output logic         [7:0]  blit_features_out, // Defines the blitter module features
    output logic         [7:0]  blit_mask_col_out, // Tells the blitter copy pixel function how to transpose the source pixel color
                                                   // Remember when writing a pixel/line/un-filled triangle/box/quad, the set color does a second
                                                   // color transpose from the copy pixel to the destination pixel color.
    output logic        [12:0]  blit_src_scale_x , // Holds the X blitter source upscale fraction, IE zoom ratio (4096:blit_src_scale_x), values 4095 through 1, or 4096 for off.
    output logic        [12:0]  blit_src_scale_y , // Holds the Y blitter source upscale fraction, IE zoom ratio (4096:blit_src_scale_y), values 4095 through 1, or 4096 for off.
    output logic        [12:0]  blit_dest_scale_x, // Holds the X blitter destination downscale fraction, IE zoom ratio (blit_dest_scale_x:4096), values 4095 through 1, or 4096 for off.
    output logic        [12:0]  blit_dest_scale_y  // Holds the Y blitter destination downscale fraction, IE zoom ratio (blit_dest_scale_y:4096), values 4095 through 1, or 4096 for off.
);

logic [1:0] sort_tri     [0:2];
logic [1:0] sort_tri_mm  [0:1];
logic [1:0] sort_quad    [0:2];
logic [1:0] sort_quad_mm [0:1];

poly_sort sorter (
// inputs
    .x_in        ( x_in      ), // values to sort
    .y_in        ( y_in      ), // values to sort
//outputs
    .sort_tri     ( sort_tri     ), // Array containing 3 sorted pointers, 1 for linegen 0 and 2 sequences for linegen 1 to generate a filled triangle using xy[0,1,2].
    .sort_tri_mm  ( sort_tri_mm  ), // Array containing 2 sorted pointers for the triangle's min Y coordinate and max Y coordinate when rendering using xy[0,1,2].
    .sort_quad    ( sort_quad    ), // Array containing 3 sorted pointers, 1 for linegen 0 and 2 sequences for linegen 1 to generate a filled triangle using xy[1,2,3].
    .sort_quad_mm ( sort_quad_mm )  // Array containing 2 sorted pointers for the triangle's min Y coordinate and max Y coordinate when rendering using xy[1,2,3].
);

logic signed [11:0] lg_out [0:3] ;  // XY output coordinates of all line generators
logic        [1:0]  lg_running   ;  // Flags stating which linegens are running
logic        [1:0]  lg_pix_rdy   ;  // Flags which linegens have ready pixels
logic        [1:0]  lg_start     ;  // Initializes the linegens to begin
logic        [1:0]  lg_pause     ;  // Freezes the lingen while they are ijn the middle of drawing
logic        [1:0]  lg_seq_cnt [0:1]  ; // Linegen sequence counters
logic        [3:0]  lg_csel    [0:3]  ; // Selects which xy[#] coordinates to use for linegen0 A,B - linegen1 A,B
logic        [3:0]  lg_csel_b  [0:3]  ; // Holds which xy[#] selection will be used for second sequence line to be drawn.

line_generator linegen_0 (
    // inputs
    .clk            ( clk                ), // 125 MHz pixel clock
    .reset          ( reset              ), // asynchronous reset
    .enable         ( enable && !blitter_busy ),  // Allows processing
    .run            ( lg_start[0]        ),       // HIGH during drawing
    .aX             ( x_in[lg_csel[2'd0][3:2]] ), // 12-bit X-coordinate for line start
    .aY             ( y_in[lg_csel[2'd0][1:0]] ), // 12-bit Y-coordinate for line start
    .bX             ( x_in[lg_csel[2'd1][3:2]] ), // 12-bit X-coordinate for line end
    .bY             ( y_in[lg_csel[2'd1][1:0]] ), // 12-bit Y-coordinate for line end
    .ena_pause      ( lg_pause[0]        ), // set HIGH to pause line generator while it is drawing
    // outputs
    .busy           ( lg_running[0]      ), // HIGH when line_generator is running
    .X_coord        ( lg_out[2'b00]      ), // 12-bit X-coordinate for current pixel
    .Y_coord        ( lg_out[2'b01]      ), // 12-bit Y-coordinate for current pixel
    .pixel_data_rdy ( lg_pix_rdy[0]      ), // HIGH when coordinate outputs are valid
    .line_complete  (                    )  // HIGH when line is completed
);

line_generator linegen_1 (
    // inputs
    .clk            ( clk                ), // 125 MHz pixel clock
    .reset          ( reset              ), // asynchronous reset
    .enable         ( enable && !blitter_busy ),  // Allows processing
    .run            ( lg_start[1]        ),       // HIGH during drawing
    .aX             ( x_in[lg_csel[2'd2][3:2]] ), // 12-bit X-coordinate for line start
    .aY             ( y_in[lg_csel[2'd2][1:0]] ), // 12-bit Y-coordinate for line start
    .bX             ( x_in[lg_csel[2'd3][3:2]] ), // 12-bit X-coordinate for line end
    .bY             ( y_in[lg_csel[2'd3][1:0]] ), // 12-bit Y-coordinate for line end
    .ena_pause      ( lg_pause[1]        ), // set HIGH to pause line generator
    // outputs
    .busy           ( lg_running[1]      ), // HIGH when line_generator is running
    .X_coord        ( lg_out[2'b10]      ), // 12-bit X-coordinate for current pixel
    .Y_coord        ( lg_out[2'b11]      ), // 12-bit Y-coordinate for current pixel
    .pixel_data_rdy ( lg_pix_rdy[1]      ), // HIGH when coordinate outputs are valid
    .line_complete  (                    )  // HIGH when line is completed
);

logic               execute_next_draw ; // goes high only when ready to accept a new command
logic               linegen_busy      ; // 
logic               fill_ena          ; // 

logic signed [11:0] y_pos             ; // Current raster Y position counter
logic signed [11:0] y_end             ; // Y raster fill ending position
logic signed [11:0] x_pos             ; // Current raster X position counter
logic signed [11:0] x_pos_bk          ; // Restore raster X position after a Y increment.
logic signed [11:0] x_end             ; // X raster fill ending coordinates
logic               rast_fill_pix_rdy ;

always_comb begin
// generate drawing processing busy flags
linegen_busy      = lg_running[0] || lg_running[1] ;
execute_next_draw = cmd_rdy_in && !blitter_busy && !plotter_busy && !fill_ena ;

// generate selection of the output write pixel port
pixel_xy[0]       = rast_fill_pix_rdy ? x_pos : (lg_out[{lg_pix_rdy[1],1'b0}]); // select between linegen0&1 X coordinates or the y_pos raster fill coordinates
pixel_xy[1]       = rast_fill_pix_rdy ? y_pos : (lg_out[{lg_pix_rdy[1],1'b1}]); // select between linegen0&1 Y coordinates or the y_pos raster fill coordinates
pixel_ena         = lg_pix_rdy[0] || lg_pix_rdy[1] || rast_fill_pix_rdy ;       // output pixel enable

end

always_ff @(posedge clk or posedge reset) begin

    if ( reset ) begin  // Reset only the key controls in the command pipe.
         blit_features_out   <= 0;
         blit_mask_col_out   <= 0;
         lg_seq_cnt[0]       <= 0;
         lg_seq_cnt[1]       <= 0;
         lg_start[0]         <= 1'b0 ;              // clear the 1-shot line start
         lg_start[1]         <= 1'b0 ;              // clear the 1-shot line start
         fill_ena            <= 1'b0 ;              // clear the 1-shot line start
         rast_fill_pix_rdy   <= 1'd0 ;
         blit_src_scale_x    <= 13'd4096 ; // Holds the X blitter source upscale fraction, 4096 = 1:1, IE disable.
         blit_src_scale_y    <= 13'd4096 ; // Holds the Y blitter source upscale fraction, 4096 = 1:1, IE disable.
         blit_dest_scale_x   <= 13'd4096 ; // Holds the X blitter destination downscale fraction, 4096 = 1:1, IE disable.
         blit_dest_scale_y   <= 13'd4096 ; // Holds the Y blitter destination downscale fraction, 4096 = 1:1, IE disable.
    end // reset
    else
    if ( enable && !blitter_busy ) begin

if (lg_start[0]) begin
  lg_seq_cnt[0] <= lg_seq_cnt[0]-1'b1; // subtract counter after linegen has been executed
  lg_start[0]   <= 1'b0 ;              // clear the 1-shot line start
  lg_csel[0]    <= lg_csel_b[0] ;      // Switch over the xy[#] selection index to the second line's coordinates
  lg_csel[1]    <= lg_csel_b[1] ;      // Switch over the xy[#] selection index to the second line's coordinates
  end
if (lg_start[1]) begin
  lg_seq_cnt[1] <= lg_seq_cnt[1]-1'b1; // subtract counter after linegen has been executed
  lg_start[1]   <= 1'b0 ;              // clear the 1-shot line start
  lg_csel[2]    <= lg_csel_b[2] ;      // Switch over the xy[#] selection index to the second line's coordinates
  lg_csel[3]    <= lg_csel_b[3] ;      // Switch over the xy[#] selection index to the second line's coordinates
  end


// ***************************************************************************************************
// Decode drawing commands and prep linegens for drawing.
// ***************************************************************************************************

if (execute_next_draw) begin
   
        if (cmd_in[15:8]  == 8'd0) blit_features_out <= cmd_in[7:0]; // Just set the blitter features
   else if (cmd_in[15:8]  == 8'd8) blit_mask_col_out <= cmd_in[7:0]; // Just set the blitter transparency mask color
   else if (cmd_in[15:8]  == 8'd9) begin                             // Set blitter scale
      if (cmd_in[0]) begin // enable setting of source scale
        if ( x_in[0]==0 )  blit_src_scale_x    <= 13'd4096        ; // If the register is 0, turn off scale factor by using 4096
        else               blit_src_scale_x    <= {1'b0,x_in[0]}  ; // Otherwize, set the scale factor to 1 through 4095.
        if ( y_in[0]==0 )  blit_src_scale_y    <= 13'd4096        ; // If the register is 0, turn off scale factor by using 4096
        else               blit_src_scale_y    <= {1'b0,y_in[0]}  ; // Otherwize, set the scale factor to 1 through 4095.
      end
      if (cmd_in[1]) begin // enable setting of source scale
        if ( x_in[1]==0 )  blit_dest_scale_x   <= 13'd4096        ; // If the register is 0, turn off scale factor by using 4096
        else               blit_dest_scale_x   <= {1'b0,x_in[1]}  ; // Otherwize, set the scale factor to 1 through 4095.
        if ( y_in[1]==0 )  blit_dest_scale_y   <= 13'd4096        ; // If the register is 0, turn off scale factor by using 4096
        else               blit_dest_scale_y   <= {1'b0,y_in[1]}  ; // Otherwize, set the scale factor to 1 through 4095.
      end
   end
   else if (cmd_in[15:12] == 4'd0) begin                             // Any other valid plotting draw command
    
        plotter_busy      <= 1 ;           // Tell the rest of the geometry processor that the plotter is going to draw
        pixel_col         <= cmd_in[7:0];  // set the output drawing color

   if ( cmd_in[10:8] == 3'd1 ) begin                 // Draw a dot
                       lg_seq_cnt[0]     <= 2'd1          ; // Linegen 0 has 1 line to draw
                       lg_csel[2'd0]     <= {2'd0,2'd0}   ; // Linegen 0's first  line's A coordinate = xy[0]
                       lg_csel[2'd1]     <= {2'd0,2'd0}   ; // Linegen 0's first  line's B coordinate = xy[0]
                       lg_csel_b[2'd0]   <= {2'd0,2'd0}   ; // Linegen 0's second line's A coordinate = xy[0]   *un-used
                       lg_csel_b[2'd1]   <= {2'd0,2'd0}   ; // Linegen 0's second line's B coordinate = xy[0]   *un-used

                       lg_seq_cnt[1]     <= 2'd0          ; // Linegen 1 has no line to draw
                       lg_csel[2'd2]     <= {2'd0,2'd0}   ; // Linegen 1's first  line's A coordinate = xy[0]   *un-used
                       lg_csel[2'd2]     <= {2'd0,2'd0}   ; // Linegen 1's first  line's B coordinate = xy[0]   *un-used
                       lg_csel_b[2'd3]   <= {2'd0,2'd0}   ; // Linegen 1's second line's A coordinate = xy[0]   *un-used
                       lg_csel_b[2'd3]   <= {2'd0,2'd0}   ; // Linegen 1's second line's B coordinate = xy[0]   *un-used

                       fill_ena          <= 1'b0   ; // turn off the filled flag

                       lg_start[0]       <= 1'b1;   // Start linegen 0 immediately.
                       lg_pause[0]       <= 1'b0;
                       lg_pause[1]       <= 1'b1;
                       end

   else if ( cmd_in[10:8] == 3'd2 ) begin                   // Draw a line
                       lg_seq_cnt[0]     <= 2'd1          ; // Linegen 0 has 1 line to draw
                       lg_csel[2'd0]     <= {2'd0,2'd0}   ; // Linegen 0's first  line's A coordinate = xy[0]
                       lg_csel[2'd1]     <= {2'd1,2'd1}   ; // Linegen 0's first  line's B coordinate = xy[1]
                       lg_csel_b[2'd0]   <= {2'd0,2'd0}   ; // Linegen 0's second line's A coordinate = xy[0]   *un-used
                       lg_csel_b[2'd1]   <= {2'd0,2'd0}   ; // Linegen 0's second line's B coordinate = xy[0]   *un-used

                       lg_seq_cnt[1]     <= 2'd0          ; // Linegen 1 has no line to draw
                       lg_csel[2'd2]     <= {2'd0,2'd0}   ; // Linegen 1's first  line's A coordinate = xy[0]   *un-used
                       lg_csel[2'd2]     <= {2'd0,2'd0}   ; // Linegen 1's first  line's B coordinate = xy[0]   *un-used
                       lg_csel_b[2'd3]   <= {2'd0,2'd0}   ; // Linegen 1's second line's A coordinate = xy[0]   *un-used
                       lg_csel_b[2'd3]   <= {2'd0,2'd0}   ; // Linegen 1's second line's B coordinate = xy[0]   *un-used

                       fill_ena          <= 1'b0   ; // turn off the filled flag
                       lg_start[0]       <= 1'b1;   // Start linegen 0 immediately.
                       lg_pause[0]       <= 1'b0;
                       lg_pause[1]       <= 1'b1;
                       end

// Vertex order of a filled triangle.
//
// xy[0]----xy[1]
//   |      /  
//   |     /       
//   |    /         
//   |   /     
//   |  /     
//   | /     
// xy[2]    xy[3] N/A
//
   else if ( cmd_in[10:8] == 3'd3 ) begin                               // Draw a triangle   *** See sorter which organizes the linegen selection
                       lg_seq_cnt[0]     <= 2'd1                      ; // Linegen 0 has 1 line to draw
                       lg_csel[2'd0]     <= {sort_tri[0],sort_tri[0]} ; // Linegen 0's first  line's A coordinate = sorted xy[0]
                       lg_csel[2'd1]     <= {sort_tri[2],sort_tri[2]} ; // Linegen 0's first  line's B coordinate = sorted xy[2]
                       lg_csel_b[2'd0]   <= {2'd0,2'd0}               ; // Linegen 0's second line's A coordinate = xy[0]   *un-used
                       lg_csel_b[2'd1]   <= {2'd0,2'd0}               ; // Linegen 0's second line's B coordinate = xy[0]   *un-used

                       lg_seq_cnt[1]     <= 2'd2                      ; // Linegen 1 has 2 lines to draw
                       lg_csel[2'd2]     <= {sort_tri[0],sort_tri[0]} ; // Linegen 1's first  line's A coordinate = sorted xy[0]
                       lg_csel[2'd3]     <= {sort_tri[1],sort_tri[1]} ; // Linegen 1's first  line's B coordinate = sorted xy[1]
                       lg_csel_b[2'd2]   <= {sort_tri[1],sort_tri[1]} ; // Linegen 1's second line's A coordinate = sorted xy[1]
                       lg_csel_b[2'd3]   <= {sort_tri[2],sort_tri[2]} ; // Linegen 1's second line's B coordinate = sorted xy[2]

                       fill_ena          <= cmd_in[11]           ; // Set the filled flag
                       y_pos             <= y_in[sort_tri_mm[0]] ; // Set the fill Y raster position starting coordinate
                       y_end             <= y_in[sort_tri_mm[1]] ; // Set the fill Y raster position ending coordinate
                       x_pos             <= x_in[sort_tri_mm[0]] ; // Set the X raster position starting coordinate
                       x_pos_bk          <= x_in[sort_tri_mm[0]] ; // Set the X raster position starting coordinate
                       x_end             <= x_in[sort_tri_mm[0]] ; // Set the X raster position ending coordinate

                       lg_start[0]       <= 1'b1;   // Start linegen 0 immediately.
                       lg_pause[0]       <= 1'b0;
                       lg_pause[1]       <= 1'b1;
                       end  // triangle

   else if ( cmd_in[10:8] == 3'd4 ) begin                 // Draw a box

// Vertex order of a non filled & filled box
//
// xy[00] -L0f- xy[10]
//   |            |       L#f means the linegen# running the first lg_csel coordinates
//  L1s          L0s
//   |            |       L#s means the linegen# running the second lg_csel_b coordinates
// xy[01] -l1f- xy[11]
//
            if (!cmd_in[11]) begin                          // A non-filled box, draw all 4 lines
                       lg_seq_cnt[0]     <= 2'd2          ; // Linegen 0 has 2 lines to draw
                       lg_csel[2'd0]     <= {2'd0,2'd0}   ; // Linegen 0's first  line's A coordinate = xy[00]
                       lg_csel[2'd1]     <= {2'd1,2'd0}   ; // Linegen 0's first  line's B coordinate = xy[10]
                       lg_csel_b[2'd0]   <= {2'd1,2'd0}   ; // Linegen 0's second line's A coordinate = xy[10]
                       lg_csel_b[2'd1]   <= {2'd1,2'd1}   ; // Linegen 0's second line's B coordinate = xy[11]

                       lg_seq_cnt[1]     <= 2'd2          ; // Linegen 1 has 2 lines to draw
                       lg_csel[2'd2]     <= {2'd1,2'd1}   ; // Linegen 1's first  line's A coordinate = xy[11]
                       lg_csel[2'd3]     <= {2'd0,2'd1}   ; // Linegen 1's first  line's B coordinate = xy[01]
                       lg_csel_b[2'd2]   <= {2'd0,2'd1}   ; // Linegen 1's second line's A coordinate = xy[01]
                       lg_csel_b[2'd3]   <= {2'd0,2'd0}   ; // Linegen 1's second line's B coordinate = xy[00]
                       end // non-filled box

// Vertex order of a filled box
//
// xy[00] **** xy[10]
//   |    ****    |
//  L0f   ****   L1f       L#f means the linegen# running the first lg_csel coordinates only
//   |    ****    |        **** is the area filled by the raster fill.
// xy[01] **** xy[11]
//
                       else begin                          // Draw the second half of a filled quadrilateral, coordinates xy[3,2,1] instead of xy[0,1,2]
                       lg_seq_cnt[0]     <= 2'd1         ; // Linegen 0 has 1 line to draw
                       lg_csel[2'd0]     <= {2'd0,2'd0}   ; // Linegen 0's first  line's A coordinate = xy[00]
                       lg_csel[2'd1]     <= {2'd0,2'd1}   ; // Linegen 0's first  line's B coordinate = xy[01]
                       lg_csel_b[2'd0]   <= {2'd0,2'd0}   ; // Linegen 0's second line's A coordinate = xy[00]   *un-used
                       lg_csel_b[2'd1]   <= {2'd0,2'd0}   ; // Linegen 0's second line's B coordinate = xy[00]   *un-used

                       lg_seq_cnt[1]     <= 2'd1          ; // Linegen 1 has 2 lines to draw
                       lg_csel[2'd2]     <= {2'd1,2'd0}   ; // Linegen 1's first  line's A coordinate = xy[10]
                       lg_csel[2'd3]     <= {2'd1,2'd1}   ; // Linegen 1's first  line's B coordinate = xy[11]
                       lg_csel_b[2'd2]   <= {2'd0,2'd0}   ; // Linegen 1's second line's A coordinate = xy[00]   *un-used
                       lg_csel_b[2'd3]   <= {2'd0,2'd0}   ; // Linegen 1's second line's B coordinate = xy[00]   *un-used
                       end  // filled box

                       fill_ena          <= cmd_in[11]  ; // Set the filled flag
                       y_pos             <= y_in[0]     ; // Set the fill Y raster position starting coordinate
                       y_end             <= y_in[1]     ; // Set the fill Y raster position ending coordinate
                       x_pos             <= x_in[0]     ; // Set the X raster position starting coordinate
                       x_pos_bk          <= x_in[0]     ; // Set the X raster position starting coordinate
                       x_end             <= x_in[1]     ; // Set the X raster position ending coordinate

                       lg_start[0]       <= 1'b1;   // Start linegen 0 immediately.
                       lg_pause[0]       <= 1'b0;
                       lg_pause[1]       <= 1'b1;
                       end // Any box

   else if ( cmd_in[10:8] == 3'd5 ) begin                 // Draw a quadrilateral

// Vertex order of a non filled quadrilateral
//
// xy[0] -L0f- xy[1]
//   |           |       L#f means the linegen# running the first lg_csel coordinates
//  L1s         L0s
//   |           |       L#s means the linegen# running the second lg_csel_b coordinates
// xy[2] -l1f- xy[3]
//
            if (!cmd_in[11]) begin                          // A non-filled quadrilateral, draw all 4 lines
                       lg_seq_cnt[0]     <= 2'd2          ; // Linegen 0 has 2 lines to draw

                       if ( y_in[0] > y_in[1] ) begin     ; // Check to see what direction line 1 of 4 would be drawn if it were drawn as a sorted quad and match it
                       lg_csel[2'd0]     <= {2'd1,2'd1}   ; // Linegen 0's first  line's A coordinate = xy[1]
                       lg_csel[2'd1]     <= {2'd0,2'd0}   ; // Linegen 0's first  line's B coordinate = xy[0]
                       end else begin                     ; // Reverse the line drawing direction for line 1 of 4.
                       lg_csel[2'd0]     <= {2'd0,2'd0}   ; // Linegen 0's first  line's A coordinate = xy[0]
                       lg_csel[2'd1]     <= {2'd1,2'd1}   ; // Linegen 0's first  line's B coordinate = xy[1]
                       end

                       if ( y_in[1] > y_in[3] ) begin     ; // Check to see what direction line 2 of 4 would be drawn if it were drawn as a sorted quad and match it
                       lg_csel_b[2'd0]   <= {2'd3,2'd3}   ; // Linegen 0's second line's A coordinate = xy[3]
                       lg_csel_b[2'd1]   <= {2'd1,2'd1}   ; // Linegen 0's second line's B coordinate = xy[1]
                       end else begin                     ; // Reverse the line drawing direction for line 2 of 4.
                       lg_csel_b[2'd0]   <= {2'd1,2'd1}   ; // Linegen 0's second line's A coordinate = xy[1]
                       lg_csel_b[2'd1]   <= {2'd3,2'd3}   ; // Linegen 0's second line's B coordinate = xy[3]
                       end

                       lg_seq_cnt[1]     <= 2'd2          ; // Linegen 1 has 2 lines to draw

                       if ( y_in[2] > y_in[3] ) begin     ; // Check to see what direction line 3 of 4 would be drawn if it were drawn as a sorted quad and match it
                       lg_csel[2'd2]     <= {2'd3,2'd3}   ; // Linegen 1's first  line's A coordinate = xy[3]
                       lg_csel[2'd3]     <= {2'd2,2'd2}   ; // Linegen 1's first  line's B coordinate = xy[2]
                       end else begin                     ; // Reverse the line drawing direction for line 3 of 4.
                       lg_csel[2'd2]     <= {2'd2,2'd2}   ; // Linegen 1's first  line's A coordinate = xy[2]
                       lg_csel[2'd3]     <= {2'd3,2'd3}   ; // Linegen 1's first  line's B coordinate = xy[3]
                       end

                       if ( y_in[0] > y_in[2] ) begin     ; // Check to see what direction line 4 of 4 would be drawn if it were drawn as a sorted quad and match it
                       lg_csel_b[2'd2]   <= {2'd2,2'd2}   ; // Linegen 1's second line's A coordinate = xy[2]
                       lg_csel_b[2'd3]   <= {2'd0,2'd0}   ; // Linegen 1's second line's B coordinate = xy[0]
                       end else begin                     ; // Reverse the line drawing direction for line 4 of 4.
                       lg_csel_b[2'd2]   <= {2'd0,2'd0}   ; // Linegen 1's second line's A coordinate = xy[0]
                       lg_csel_b[2'd3]   <= {2'd2,2'd2}   ; // Linegen 1's second line's B coordinate = xy[2]
                       end

                       end // non-filled quadrilateral

// Vertex order of a filled quadrilateral, command sent after filled triangle.
// *** xy[0,1,2] was drawn with a filled triangle
//
// xy[0]    xy[1]
//  N/A     / |
//         /  |    *** See sorter which organizes the linegen selection
//        /   |        Subtract 1 for each position
//       /    |
// xy[2] -- xy[3]
//
                       else begin                                         // Draw the second half of a filled quadrilateral, coordinates xy[1,2,3] instead of xy[0,1,2]
                       lg_seq_cnt[0]     <= 2'd1                        ; // Linegen 0 has 1 line to draw
                       lg_csel[2'd0]     <= {sort_quad[0],sort_quad[0]} ; // Linegen 0's first  line's A coordinate = sorted xy[0]
                       lg_csel[2'd1]     <= {sort_quad[2],sort_quad[2]} ; // Linegen 0's first  line's B coordinate = sorted xy[2]
                       lg_csel_b[2'd0]   <= {2'd0,2'd0}                 ; // Linegen 0's second line's A coordinate = xy[0]   *un-used
                       lg_csel_b[2'd1]   <= {2'd0,2'd0}                 ; // Linegen 0's second line's B coordinate = xy[0]   *un-used

                       lg_seq_cnt[1]     <= 2'd2                        ; // Linegen 1 has 2 lines to draw
                       lg_csel[2'd2]     <= {sort_quad[0],sort_quad[0]} ; // Linegen 1's first  line's A coordinate = sorted xy[0]
                       lg_csel[2'd3]     <= {sort_quad[1],sort_quad[1]} ; // Linegen 1's first  line's B coordinate = sorted xy[1]
                       lg_csel_b[2'd2]   <= {sort_quad[1],sort_quad[1]} ; // Linegen 1's second line's A coordinate = sorted xy[1]
                       lg_csel_b[2'd3]   <= {sort_quad[2],sort_quad[2]} ; // Linegen 1's second line's B coordinate = sorted xy[2]
                       end  // filled quadrilateral

                       fill_ena          <= cmd_in[11]            ; // Set the filled flag
                       y_pos             <= y_in[sort_quad_mm[0]] ; // Set the Y raster position starting coordinate
                       y_end             <= y_in[sort_quad_mm[1]] ; // Set the Y raster position ending coordinate
                       x_pos             <= x_in[sort_quad_mm[0]] ; // Set the X raster position starting coordinate
                       x_pos_bk          <= x_in[sort_quad_mm[0]] ; // Set the X raster position starting coordinate
                       x_end             <= x_in[sort_quad_mm[0]] ; // Set the X raster position ending coordinate

                       lg_start[0]       <= 1'b1;   // Start linegen 0 immediately.
                       lg_pause[0]       <= 1'b0;
                       lg_pause[1]       <= 1'b1;
                       end // Any Quadrilateral

   end // Any other valid plotting draw command
end // if (execute_next_draw)

   else if (plotter_busy) begin // A draw plot command is to be run

  if ( !fill_ena  ) begin // run the 2 linegens in a sequential manner, 1 after the other.

if (!linegen_busy) begin
      if ( lg_seq_cnt[0]!=0 ) begin      // If there are sequences, first run linegen 0
      lg_start[0]   <= 1'b1;
      lg_pause[0]   <= 1'b0;
      lg_pause[1]   <= 1'b1;
      end 
      else if ( lg_seq_cnt[1]!=0 ) begin // Then, if there are sequences for linegen 1, cycle them.
      lg_start[1]   <= 1'b1;
      lg_pause[0]   <= 1'b1;
      lg_pause[1]   <= 1'b0;
      end
       // Nothing left to draw, so, exit plotter_busy
       else if (!linegen_busy && lg_seq_cnt[0]==0 && lg_seq_cnt[1]==0 ) plotter_busy  <= 0 ;
    end
       // If linegen1 is finished and linegen0 isn't but it is paused, un-pause it.
       else if (!lg_running[1] && lg_seq_cnt[1]==0 && lg_running[0] && lg_pause[0] ) lg_pause[0] <= 0;
       // If linegen0 is finished and linegen1 isn't but it is paused, un-pause it.
       else if (!lg_running[0] && lg_seq_cnt[0]==0 && lg_running[1] && lg_pause[1] ) lg_pause[1] <= 0;

   end else begin // run the 2 linegens in a parallel fashion aligning them to a Y raster counter & fill a horizontal line between the X coordinates

if (fill_ena)
   if (!lg_running[0] && lg_seq_cnt[0]!=0 && !lg_start[1] && !lg_pause[0]) begin
         lg_start[0]       <= 1'b1;
         lg_pause[0]       <= 1'b0;
         lg_pause[1]       <= 1'b1;
   end else if (!lg_running[1] && lg_seq_cnt[1]!=0 && !lg_start[0] && !lg_pause[1]) begin
         lg_start[1]       <= 1'b1;
         lg_pause[0]       <= 1'b1;
         lg_pause[1]       <= 1'b0;
   end else begin

    if (lg_pause==2'd3) begin                              // If both linegens as paused simultaneously because both of their output Y coordinates
                                                           // sent a coordinate matching the current raster fill coordinate y_pos.
         
          if (x_pos != x_end) begin                        // if there is a void in-between the 2 linegen's X coordinates
               rast_fill_pix_rdy <= 1'b1;                  // Switch output draw pixel coordinates from linegens to fill x&y_pos coordinates
               if (x_pos > x_end ) x_pos <= x_pos - 1'b1;  // inc/dec X fill coordinate.
               else                x_pos <= x_pos + 1'b1;

           end else begin                               // if the fill is finished or there was nothing to fill

           rast_fill_pix_rdy <= 1'b0;                   // Switch output draw pixel coordinates from raster fill x&y_pos back to linegen outputs.

           if (y_pos == y_end) fill_ena <= 1'b0 ;       // if we have filled the last line, then end the flodd fill.

               if (y_pos > y_end ) y_pos <= y_pos - 1'b1;  // inc/dec X fill coordinate.
               else                y_pos <= y_pos + 1'b1;
                                   x_pos <= x_pos_bk ;     // restore X position after Y increment.

           if (lg_running[0] || lg_seq_cnt[0]!=0) lg_pause <= 2'd2; // if linegen 0 still has work to do, re-start linegen 0, freeze linegen 1
           else                                   lg_pause <= 2'd1; // Otherwise, continue linegen 1 if it has any remaining pixels.
           
           end

    end else begin

           if (lg_out[2'b01][1:0] == y_pos[1:0] && lg_pix_rdy[0] ) begin        // if linegen 0 outputs a valid Y coordinate matching the y_pos[0]
                                                 lg_pause[0] <= 1'b1;           // pause linegen 0
                                                 lg_pause[1] <= 1'b0;           // un-pause linegen 1
                                                 x_pos       <= lg_out[2'b00] ; // set the initial X fill coordinate counter
                                                 x_pos_bk    <= lg_out[2'b00] ; // set the initial X fill coordinate counter backup return position
                                                 end

           if (lg_out[2'b11][1:0] == y_pos[1:0] && lg_pix_rdy[1] ) begin        // if linegen 1 outputs a valid Y coordinate matching the y_pos[0]
                                                 lg_pause[1] <= 1'b1;           // pause linegen 1
                                                 
                                                 // This trick eliminates the linegen1's last written pixel from the raster fill by incrementing the x_end position once in the
                                                 // correct direction only if needed before the fill algorithm begins which checks to see if x_pos & x_end are equal before beginning
                                                          if (x_pos_bk == lg_out[2'b10] ) x_end       <= lg_out[2'b10]       ;  // Keep equal coordinate
                                                     else if (x_pos_bk <  lg_out[2'b10] ) x_end       <= lg_out[2'b10] - 1'b1;  // inc/dec X fill final coordinate.
                                                     else                                 x_end       <= lg_out[2'b10] + 1'b1;
                                                 end

         end
         
   end
   
end
   
   end // plotter busy loop
 end // enable
end // always_ff

endmodule



/*
 * poly_sort module
 *
 * Outputs pointer which control the selection of xy[#'s]
 * each linegen 0&1 will use to draf a filled tri and filled quad
 * Also outputs pointers to the min and max Y coords in
 * the filled triangle and filled quad
 *
 */

module poly_sort (
// inputs
    input  logic signed [11:0] x_in [0:3]         , // values to sort
    input  logic signed [11:0] y_in [0:3]         , // values to sort
//outputs
    output logic        [1:0]  sort_tri     [0:2] , // Array containing 3 sorted pointers, 1 for linegen 0 and 2 sequences for linegen 1 to generate a filled triangle using xy[0,1,2].
    output logic        [1:0]  sort_tri_mm  [0:1] , // Array containing 2 sorted pointers for the triangle's min Y coordinate and max Y coordinate when rendering using xy[0,1,2].
    output logic        [1:0]  sort_quad    [0:2] , // Array containing 3 sorted pointers, 1 for linegen 0 and 2 sequences for linegen 1 to generate a filled triangle using xy[1,2,3].
    output logic        [1:0]  sort_quad_mm [0:1]   // Array containing 2 sorted pointers for the triangle's min Y coordinate and max Y coordinate when rendering using xy[3,2,1].
);

always_comb begin

// *********************************************************************
// Copy the Y sort to the correct line generators for a filled triangle
// *********************************************************************
//   xy[0]
//    ***
//    *  LG1f        f = first of 2 lines to draw
//    *    ** 
//   LG0f   xy[1]
//    *    **
//    *  LG1s        s = second of 2 lines to draw
//    ***
//   xy[2]           LG0 only draws 1 line
//
sort_tri_mm[1'b0] = sort_tri[0] ; // Triangle minimum Y coordinate
sort_tri_mm[1'b1] = sort_tri[2] ; // Triangle minimum Y coordinate

// *********************************************************************
// Copy the Y sort to the correct line generators for a filled quad
// *********************************************************************
//   xy[1]
//    ***
//    *  LG1f        f = first of 2 lines to draw
//    *    ** 
//   LG0f   xy[2]
//    *    **
//    *  LG1s        s = second of 2 lines to draw
//    ***
//   xy[3]           LG0 only draws 1 line
//
sort_quad_mm[1'b0] = sort_quad[0] ; // Quad minimum Y coordinate
sort_quad_mm[1'b1] = sort_quad[2] ; // Quad minimum Y coordinate

// ***************************************************
// Generate the Y order for the sorted triangle
// ***************************************************

            if ( ( y_in[0] >=  y_in[1] ) && ( y_in[1] >= y_in[2] ) ) begin
                sort_tri[0] = 2'd2 ;
                sort_tri[1] = 2'd1 ;
                sort_tri[2] = 2'd0 ;
            end else
            if ( ( y_in[1] >=  y_in[2] ) && ( y_in[2] >= y_in[0] ) ) begin
                sort_tri[0] = 2'd0 ;
                sort_tri[1] = 2'd2 ;
                sort_tri[2] = 2'd1 ;
            end else
            if ( ( y_in[2] >=  y_in[0] ) && ( y_in[0] >= y_in[1] ) ) begin
                sort_tri[0] = 2'd1 ;
                sort_tri[1] = 2'd0 ;
                sort_tri[2] = 2'd2 ;
            end else
            if ( ( y_in[0] >=  y_in[2] ) && ( y_in[2] >= y_in[1] ) ) begin
                sort_tri[0] = 2'd1 ;
                sort_tri[1] = 2'd2 ;
                sort_tri[2] = 2'd0 ;
            end else
            if ( ( y_in[2] >=  y_in[1] ) && ( y_in[1] >= y_in[0] ) ) begin
                sort_tri[0] = 2'd0 ;
                sort_tri[1] = 2'd1 ;
                sort_tri[2] = 2'd2 ;
            end else
            if ( ( y_in[1] >=  y_in[0] ) && ( y_in[0] >= y_in[2] ) ) begin
                sort_tri[0] = 2'd2 ;
                sort_tri[1] = 2'd0 ;
                sort_tri[2] = 2'd1 ;
            end
// ***************************************************        
// Generate the Y order for the sorted quad
// *************************************************** 
       
            if ( ( y_in[1] >=  y_in[2] ) && ( y_in[2] >= y_in[3] ) ) begin
                sort_quad[0] = 2'd3 ;
                sort_quad[1] = 2'd2 ;
                sort_quad[2] = 2'd1 ;
            end else
            if ( ( y_in[2] >=  y_in[3] ) && ( y_in[3] >= y_in[1] ) ) begin
                sort_quad[0] = 2'd1 ;
                sort_quad[1] = 2'd3 ;
                sort_quad[2] = 2'd2 ;
            end else
            if ( ( y_in[3] >=  y_in[1] ) && ( y_in[1] >= y_in[2] ) ) begin
                sort_quad[0] = 2'd2 ;
                sort_quad[1] = 2'd1 ;
                sort_quad[2] = 2'd3 ;
            end else
            if ( ( y_in[1] >=  y_in[3] ) && ( y_in[3] >= y_in[2] ) ) begin
                sort_quad[0] = 2'd2 ;
                sort_quad[1] = 2'd3 ;
                sort_quad[2] = 2'd1 ;
            end else
            if ( ( y_in[3] >=  y_in[2] ) && ( y_in[2] >= y_in[1] ) ) begin
                sort_quad[0] = 2'd1 ;
                sort_quad[1] = 2'd2 ;
                sort_quad[2] = 2'd3 ;
            end else
            if ( ( y_in[2] >=  y_in[1] ) && ( y_in[1] >= y_in[3] ) ) begin
                sort_quad[0] = 2'd3 ;
                sort_quad[1] = 2'd1 ;
                sort_quad[2] = 2'd2 ;
            end

end
=======
                    draw_cmd_func        <= CMD_OUT_RST_PXWRI_M[3:0];                   // sets the output funtion
                    draw_cmd_data_color  <= command_data8;                              // sets the mask color
                    draw_cmd_data_word_Y <= { command_data8[7:0], command_data8[7:4] }; // sets mask color #2 and 1/2 or #3
                    draw_cmd_data_word_X <= { command_data8[3:0], command_data8[7:4] }; // sets mask color 1/2 or #3 and #4
                    draw_cmd_tx          <= 1'b1;                                       // transmits the command
                end
                
                8'd90 : begin               // clear the blitter copy pixel collision counter
                    draw_cmd_func        <= CMD_OUT_RST_PXPASTE_M[3:0];                 // sets the output funtion
                    draw_cmd_data_color  <= command_data8;                              // sets the mask color
                    draw_cmd_data_word_Y <= { command_data8[7:0], command_data8[7:4] }; // sets mask color #2 and 1/2 or #3
                    draw_cmd_data_word_X <= { command_data8[3:0], command_data8[7:4] }; // sets mask color 1/2 or #3 and #4
                    draw_cmd_tx          <= 1'b1;                                       // transmits the command
                end

                8'b000????? : begin // this range of commands all begin drawing a shape
                
               // drawing commands begin here.  Keep the convention that:
               // extend_cmd[3] = fill enable
               // extend_cmd[4] = use the color in the copy/paste buffer.  This one is for drawing in true color mode.
               // extend_cmd[5] = mask enable - when drawing, the mask colours will not be plotted as they are transparent
                    geo_shape[3]         <= 1'b0;               // geo shapes 0 through 7, geo shapes 8 through 15 are for copy & paste.
                    geo_shape[2:0]       <= command_in[2:0];    // Set which one of shapes 0 through 7 should be drawn.  Shape 0 means nothing is being drawn
                    geo_fill             <= command_in[3];      // Fill enable bit
                    geo_paste            <= command_in[4];      // Used for drawing in true color 16 bit mode
                    geo_mask             <= 1'b0;               // Mask disables when drawing raw geometry shapes
                    geo_run              <= 1'b1;               // A flag which signifies that a geometric shape drawing engine will begin drawing
                    geo_color            <= command_data8;      // set the 8-bit pen color
                    
                    if ( command_in[2:0] == 4'd1 ) linegen_start <= 1'b1 ;  // Start line_generator to draw a line
                    
                    geo_sub_func1        <= 4'b0;               // for geometric engines which have multiple phases, reset the phase counter
                    geo_sub_func2        <= 4'b0;               // for geometric engines which have 2-dimensional multiple phases, reset the phase counter
                    
                    // Initialize the geometry unit starting coordinates and direction so it can begin plotting immediately
                    geo_x                <= x[0];               // initialize the beginning pixel location
                    geo_y                <= y[0];               // initialize the beginning pixel location
                    if ( x[1] < x[0] ) geo_xdir <= 12'd0-12'd1; // set the direction of the counter (negative x in this case)
                    else if ( x[1] == x[0]) geo_xdir <= 12'd0;  // neutral x direction
                    else               geo_xdir <= 12'd1;       // positive x direction
                    if ( y[1] < y[0] ) geo_ydir <= 12'd0-12'd1; // negative y direction
                    else if ( y[1] == y[0]) geo_ydir <= 12'd0;  // neutral y direction
                    else               geo_ydir <= 12'd1;       // positive y direction
                    
                    dx <= (x[1]>x[0]) ? (x[1]-x[0]) : (x[0]-x[1]); // get absolute size of delta-x
                    dy <= (y[0]>y[1]) ? (y[1]-y[0]) : (y[0]-y[1]); // get absolute size of delta-y
                    
                end

                default : begin
                
                    draw_cmd_tx <= 1'b0 ; // stop transmit output command function
                    geo_shape   <= 4'b0 ; // turn off the drawing shape
                    
                end
                
            endcase
            
        end else if ( geo_run ) begin

            case (geo_shape)    // run a selected geometric drawing engine

                4'd1 : begin    // draw line from (x[0],y[0]) to (x[1],y[1])
                        
				   draw_cmd_func        <= CMD_OUT_PXWRI[3:0] ;// Set up command to pixel plotter to write a pixel,
				   draw_cmd_data_color  <= geo_color ;         // ... in geo_colour,
				   pass_thru_a          <= 1'b0  ;
				   pass_thru_b          <= 1'b0  ;
				   draw_cmd_data_word_Y <= gen_y ;             // ... at Y-coordinate,
				   draw_cmd_data_word_X <= gen_x ;             // ... and X-coordinate.

				   if ( line_dat_rdy && ( draw_cmd_data_word_X >= 0 && draw_cmd_data_word_X <= max_x ) && ( draw_cmd_data_word_Y >=0 && draw_cmd_data_word_X <= max_y ) )
					  draw_cmd_tx       <= 1'b1  ;             // send command if geo_X&Y are within valid drawing area
				   else
					  draw_cmd_tx       <= 1'b0  ;             // otherwise turn off draw command
				   
				   if ( line_done ) begin
				   
					  geo_shape     <= 4'd0 ; // last pixel
					  linegen_start <= 1'b0 ; // reset linegen_start
					  
				   end
                
                end // geo_shape - draw line
                
                4'd2 : begin    // draw a filled rectangle

                    if ( geo_y != (y[1] + geo_ydir) ) begin              // Check for bottom (or top, depending on sign of geo_ydir) of rectangle reached
                    
                        if ( geo_x != (x[1] + geo_xdir) ) begin          // Check for right (or left, depending on sign of geo_xdir) of rectangle reached
                        
                            draw_cmd_func        <= CMD_OUT_PXWRI[3:0] ; // Set up command to pixel plotter to write a pixel,
                            draw_cmd_data_color  <= geo_color ;          // ... in geo_colour,
                            draw_cmd_data_word_Y <= geo_y     ;          // ... at Y-coordinate,
                            draw_cmd_data_word_X <= geo_x     ;          // ... and X-coordinate.
                            
                            if ( (geo_x >= 0 && geo_x <= max_x) && (geo_y >= 0 && geo_y <= max_y) )
                                draw_cmd_tx  <= 1'b1 ; // send command if geo_X&Y are within valid drawing area
                            else
                                draw_cmd_tx  <= 1'b0 ; // otherwise turn off draw command
                            
                            // Now increment (or decrement according to geo_xdir) geo_x to the next pixel.
                            // If geo_fill is HIGH, step to next X-position to fill the rectangle.
                            // If geo_x is at the end edge, step past it.
                            // If geo_y is at start or end (top or bottom edge), step to next X-position to draw the horizontal line.
                            if (geo_fill || geo_x == x[1] || geo_y == y[0] || geo_y == y[1] )   geo_x <= geo_x + geo_xdir ;
                            // Otherwise, jump to end X-position to draw other edge for non-filled rectangle.
                            else                                                                geo_x <= x[1] ;

                        end else begin  // geo_x has passed vertical edge
                        
                            draw_cmd_tx         <= 1'b0 ;               // do not send a draw cmd this cycle
                            geo_x               <= x[0] ;               // reset X to start X-position
                            geo_y               <= geo_y + geo_ydir ;   // increment (or decrement) Y-position for next line
                            
                        end
                    end else begin      // geo_y has passed horizontal edge
                    
                            geo_run             <= 1'b0 ;               // stop geometry engine - shape completed
                            draw_cmd_tx         <= 1'b0 ;               // do not send a draw cmd this cycle
                            
                    end
                    
                end // draw a filled rectangle

                default : begin
                
                    geo_run         <= 1'b0 ; // no valid drawing engine selected, so stop the geo_run flag.
                    draw_cmd_tx     <= 1'b0 ;
                    
                end

            endcase   // run a selected geometric drawing engine
                
        end else   draw_cmd_tx <= 1'b0 ;    // stop transmit output command function//  end of (geo_run) flag
    
    end // !draw_busy

end //always @(posedge clk)

endmodule

module tri_comp (

// inputs
   input  logic                    clk,
   input  logic signed [3:0][11:0] in,
// outputs
   output logic        [15:0]      in_a_eq_b,
   output logic        [15:0]      in_a_gt_b,
   output logic        [15:0]      in_a_lt_b

);

parameter bit CLOCK_OUTPUT = 0;

always_comb begin

   if ( ~CLOCK_OUTPUT ) begin
   
      for (int i = 0 ; i<=15 ; i++) begin
      
         in_a_eq_b[i] = ( in[ i[3:2] ] == in[ i[1:0] ] ) ;
         in_a_gt_b[i] = ( in[ i[3:2] ] >  in[ i[1:0] ] ) ;
         in_a_lt_b[i] = ( in[ i[3:2] ] <  in[ i[1:0] ] ) ;
         
      end
      
   end

end

always_ff @( posedge clk ) begin

   if ( CLOCK_OUTPUT ) begin
   
      for (int i = 0 ; i<=15 ; i++) begin
      
         in_a_eq_b[i] <= ( in[ i[3:2] ] == in[ i[1:0] ] ) ;
         in_a_gt_b[i] <= ( in[ i[3:2] ] >  in[ i[1:0] ] ) ;
         in_a_lt_b[i] <= ( in[ i[3:2] ] <  in[ i[1:0] ] ) ;
         
      end
      
   end

end

>>>>>>> e95a3e278b115b0ea9f980c63d48b6bfbcc232d1
endmodule
