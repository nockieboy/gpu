// *** Table begin.

localparam int dlut_8  [0:31] = '{     0,     1,     2,     3,     4,     5,     6,     8,    10,    12,    14,    17,    19,    23,    26,    31,    35,    41,    47,    54,    62,    70,    80,    92,   104,   119,   135,   154,   175,   198,   225,   255};
localparam int dlut_9  [0:31] = '{     0,     1,     2,     3,     4,     6,     8,    10,    13,    15,    19,    22,    27,    32,    38,    45,    53,    62,    72,    84,    99,   115,   134,   156,   181,   210,   244,   283,   328,   381,   441,   511};
localparam int dlut_10 [0:31] = '{     0,     1,     2,     4,     5,     7,    10,    13,    16,    20,    25,    30,    37,    44,    54,    64,    77,    92,   110,   132,   157,   186,   221,   263,   312,   370,   439,   520,   616,   730,   864,  1023};
localparam int dlut_11 [0:31] = '{     0,     1,     3,     4,     6,     9,    12,    16,    20,    26,    32,    40,    50,    61,    75,    92,   113,   137,   167,   204,   248,   301,   365,   442,   536,   650,   787,   953,  1154,  1397,  1691,  2047};
localparam int dlut_12 [0:31] = '{     0,     1,     3,     5,     8,    11,    15,    19,    25,    33,    42,    53,    67,    84,   105,   131,   163,   203,   253,   314,   390,   484,   600,   743,   920,  1140,  1411,  1746,  2161,  2675,  3310,  4095};
localparam int dlut_13 [0:31] = '{     0,     1,     3,     6,     9,    13,    17,    24,    31,    41,    53,    69,    89,   114,   145,   185,   236,   300,   381,   483,   613,   776,   983,  1245,  1577,  1996,  2526,  3197,  4045,  5118,  6475,  8191};
localparam int dlut_14 [0:31] = '{     0,     2,     4,     7,    10,    15,    21,    28,    38,    51,    68,    90,   118,   154,   201,   261,   340,   441,   572,   742,   961,  1245,  1612,  2086,  2700,  3494,  4521,  5849,  7568,  9790, 12665, 16383};

localparam int dlut_sel [8:14][0:31] = '{ dlut_8, dlut_9, dlut_10, dlut_11, dlut_12, dlut_13, dlut_14 };

// *** Table End.

